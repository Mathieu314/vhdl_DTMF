0
3
6
9
12
15
17
20
22
24
26
27
29
30
30
31
31
31
30
30
29
27
26
24
22
20
17
15
12
9
6
3
0
-3
-6
-9
-12
-15
-17
-20
-22
-24
-26
-27
-29
-30
-30
-31
-31
-31
-30
-30
-29
-27
-26
-24
-22
-20
-17
-15
-12
-9
-6
-3
